grammar edu:umn:cs:melt:exts:ableC:prolog;

{--
 - Here we export the concrete and abstract syntax of this extension in the
 - top-level extension grammar, so that an extension user can simply add this
 - grammar to a parser specification, or an extension writer can import both the
 - abstract syntax and concrete syntax of an extension by importing this grammar.
 -}
exports edu:umn:cs:melt:exts:ableC:prolog:core;
exports edu:umn:cs:melt:exts:ableC:prolog:list;

