grammar edu:umn:cs:melt:exts:ableC:prolog:core;

exports edu:umn:cs:melt:exts:ableC:prolog:core:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:prolog:core:concretesyntax;

