grammar edu:umn:cs:melt:exts:ableC:prolog:list;

exports edu:umn:cs:melt:exts:ableC:prolog:list:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:prolog:list:concretesyntax;

